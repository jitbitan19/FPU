`timescale 1ns / 1ps

module fp_div(a, b, ra, q, qFlags, exception);

  
endmodule