module fp_class (
    nan, inf, zero, dnorm, norm // output
    f // input
);
    parameter nexp = 11;
    parameter nman = 52;
    parameter bias = 1<<(nexp-1);
    


    input
    
endmodule